-------------------------------------------------------------------------------
--
-- Title       : R3_instruction
-- Design      : MIPS
-- Author      : Dongyun Lee
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : //Mac/Home/Documents/SBU_2024_Fall/ESE345/ese345_project/ese345_project/MIPS/src/R3_instruction.vhd
-- Generated   : Mon Oct 21 16:29:10 2024
-- From        : Interface description file
-- By          : ItfToHdl ver. 1.0
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--    and may be overwritten
--{entity {R3_instruction} architecture {R3_instruction}}



entity R3_instruction is
end R3_instruction;

--}} End of automatically maintained section

architecture R3_instruction of R3_instruction is
begin

	-- Enter your statements here --

end R3_instruction;
